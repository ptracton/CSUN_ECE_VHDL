-------------------------------------------------------------------------------
-- Title      : Zybo Z7010 Board Package
-- Project    : 
-------------------------------------------------------------------------------
-- File       : zybo_pkg.vhd
-- Author     : Phil Tracton  <ptracton@gmail.com>
-- Company    : CSUN
-- Created    : 2023-08-31
-- Last update: 2023-09-01
-- Platform   : Modelsim on Linux
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2023 CSUN
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2023-08-31  1.0      ptracton	Created
-------------------------------------------------------------------------------

package board_pkg is

  -- This is for the Arty S7 which has 4 switches and LEDs
  constant WIDTH : integer := 4;
  
end package;

