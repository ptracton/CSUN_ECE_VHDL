-------------------------------------------------------------------------------
-- Title      : Boolean Board GPIO
-- Project    : 
-------------------------------------------------------------------------------
-- File       : boolean_pkg.vhd
-- Author     : Phil Tracton  <ptracton@gmail.com>
-- Company    : 
-- Created    : 2025-03-05
-- Last update: 2025-03-05
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: 
-------------------------------------------------------------------------------
-- Copyright (c) 2025 
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Version  Author  Description
-- 2025-03-05  1.0      ptracton	Created
-------------------------------------------------------------------------------

package board_pkg is

  -- This is for the boolean board which has 16 Switches and LEDs
  constant WIDTH : integer := 16;
  
end package;
